-------------------------------------------------------------------------------
--
-- Title       : pseudorng
-- Design      : pseudorng_design
-- Author      : 
-- Company     : 
--
-------------------------------------------------------------------------------
--
-- File        : pseudorng.vhd
-- Generated   : Thu May 17 21:34:17 2018
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {pseudorng} architecture {asdas}}

library IEEE;
use IEEE.STD_LOGIC_1164.all;
